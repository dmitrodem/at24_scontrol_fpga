`default_nettype none
module pll (
  input wire clkin,
  input wire reset,
  output wire clkout,
  output wire locked
);
  wire gnd;
  assign gnd = 1'b0;
  PLLA #(
    // Parameters
    .FCLKIN                        ("50"),
    .IDIV_SEL                      (1),
    .FBDIV_SEL                     (1),
    .ODIV0_SEL                     (14),
    .ODIV1_SEL                     (8),
    .ODIV2_SEL                     (8),
    .ODIV3_SEL                     (8),
    .ODIV4_SEL                     (8),
    .ODIV5_SEL                     (8),
    .ODIV6_SEL                     (8),
    .MDIV_SEL                      (14),
    .MDIV_FRAC_SEL                 (0),
    .ODIV0_FRAC_SEL                (0),
    .CLKOUT0_EN                    ("TRUE"),
    .CLKOUT1_EN                    ("FALSE"),
    .CLKOUT2_EN                    ("FALSE"),
    .CLKOUT3_EN                    ("FALSE"),
    .CLKOUT4_EN                    ("FALSE"),
    .CLKOUT5_EN                    ("FALSE"),
    .CLKOUT6_EN                    ("FALSE"),
    .CLKFB_SEL                     ("INTERNAL"),
    .CLKOUT0_DT_DIR                (1'b1),
    .CLKOUT1_DT_DIR                (1'b1),
    .CLKOUT2_DT_DIR                (1'b1),
    .CLKOUT3_DT_DIR                (1'b1),
    .CLKOUT0_DT_STEP               (1'b0),
    .CLKOUT1_DT_STEP               (1'b0),
    .CLKOUT2_DT_STEP               (1'b0),
    .CLKOUT3_DT_STEP               (1'b0),
    .CLK0_IN_SEL                   (1'b0),
    .CLK0_OUT_SEL                  (1'b0),
    .CLK1_IN_SEL                   (1'b0),
    .CLK1_OUT_SEL                  (1'b0),
    .CLK2_IN_SEL                   (1'b0),
    .CLK2_OUT_SEL                  (1'b0),
    .CLK3_IN_SEL                   (1'b0),
    .CLK3_OUT_SEL                  (1'b0),
    .CLK4_IN_SEL                   (1'b0),
    .CLK4_OUT_SEL                  (1'b0),
    .CLK5_IN_SEL                   (1'b0),
    .CLK5_OUT_SEL                  (1'b0),
    .CLK6_IN_SEL                   (1'b0),
    .CLK6_OUT_SEL                  (1'b0),
    .DYN_DPA_EN                    ("FALSE"),
    .CLKOUT0_PE_COARSE             (0),
    .CLKOUT0_PE_FINE               (0),
    .CLKOUT1_PE_COARSE             (0),
    .CLKOUT1_PE_FINE               (0),
    .CLKOUT2_PE_COARSE             (0),
    .CLKOUT2_PE_FINE               (0),
    .CLKOUT3_PE_COARSE             (0),
    .CLKOUT3_PE_FINE               (0),
    .CLKOUT4_PE_COARSE             (0),
    .CLKOUT4_PE_FINE               (0),
    .CLKOUT5_PE_COARSE             (0),
    .CLKOUT5_PE_FINE               (0),
    .CLKOUT6_PE_COARSE             (0),
    .CLKOUT6_PE_FINE               (0),
    .DYN_PE0_SEL                   ("FALSE"),
    .DYN_PE1_SEL                   ("FALSE"),
    .DYN_PE2_SEL                   ("FALSE"),
    .DYN_PE3_SEL                   ("FALSE"),
    .DYN_PE4_SEL                   ("FALSE"),
    .DYN_PE5_SEL                   ("FALSE"),
    .DYN_PE6_SEL                   ("FALSE"),
    .DE0_EN                        ("FALSE"),
    .DE1_EN                        ("FALSE"),
    .DE2_EN                        ("FALSE"),
    .DE3_EN                        ("FALSE"),
    .DE4_EN                        ("FALSE"),
    .DE5_EN                        ("FALSE"),
    .DE6_EN                        ("FALSE"),
    .RESET_I_EN                    ("FALSE"),
    .RESET_O_EN                    ("FALSE"),
    .ICP_SEL                       (6'bxxxxxx),
    .LPF_RES                       (3'bxxx),
    .LPF_CAP                       (2'b00),
    .SSC_EN                        ("FALSE"))
  u0 (/*AUTOINST*/
    // Outputs
    .MDRDO            (),
    .LOCK             (locked),
    .CLKOUT0          (clkout),
    .CLKOUT1          (),
    .CLKOUT2          (),
    .CLKOUT3          (),
    .CLKOUT4          (),
    .CLKOUT5          (),
    .CLKOUT6          (),
    .CLKFBOUT         (),
    // Inputs
    .CLKIN            (clkin),
    .CLKFB            (gnd),
    .RESET            (reset),
    .PLLPWD           (gnd),
    .RESET_I          (gnd),
    .RESET_O          (gnd),
    .PSSEL            ({gnd, gnd, gnd}),
    .PSDIR            (gnd),
    .PSPULSE          (gnd),
    .SSCPOL           (gnd),
    .SSCON            (gnd),
    .SSCMDSEL         ({gnd, gnd, gnd, gnd, gnd, gnd, gnd}),
    .SSCMDSEL_FRAC    ({gnd, gnd, gnd}),
    .MDCLK            (gnd),
    .MDOPC            ({gnd, gnd}),
    .MDAINC           (gnd),
    .MDWDI            ({gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd}));
endmodule
`default_nettype wire

// Local Variables:
// verilog-library-directories: ("." "src")
// End:
